module main (output v6c86ce);
 wire w0;
 assign v6c86ce = w0;
 main_bit_1 vd05a21 (
  .v608bd9(w0)
 );
endmodule

module main_bit_1 (output v608bd9);
 wire w0;
 assign v608bd9 = w0;
 main_bit_1_basic_code_v68c173 v68c173 (
  .v(w0)
 );
endmodule

module main_bit_1_basic_code_v68c173 (output v);
 // Bit 1
 
 assign v = 1'b1;
endmodule

